`timescale 1ns / 1ps
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Company:    Penn State    	
//					
// Engineer: Marc Khouri & Matt Henry
//
// Create Date:	3/23/14
// Design Name: register_file.v
// Module Name: register_file
// Project Name: MIPS CPU
//
// Dependencies:
//
// Revision: 1
//
//
// Additional Comments:
//
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module register_file
(
    //--------------------------
	// Input Ports
	//--------------------------
	input					clk,
    input 		[4:0]		raddr0,
	input 		[4:0]		raddr1,
	input 		[4:0]		waddr,
	input		[31:0]		wdata,
	input 					wren,
    //--------------------------
    // Output Ports
    //--------------------------
    output 		[31:0] 		rdata0,
	output		[31:0]		rdata1
);
      
    ///////////////////////////////////////////////////////////////////
    // Begin Design
    ///////////////////////////////////////////////////////////////////
    //-------------------------------------------------
    // Signal Declarations: local params
    //-------------------------------------------------
	
    //-------------------------------------------------
    // Signal Declarations: reg
    //-------------------------------------------------
	reg [31:0] register_file[0:31];
	
    //-------------------------------------------------
    // Signal Declarations: wire
    //-------------------------------------------------
		
	//---------------------------------------------------------------
	// Instantiations
	//---------------------------------------------------------------
	// None

	//---------------------------------------------------------------
	// Combinatorial Logic
	//---------------------------------------------------------------

	assign rdata0 = register_file[raddr0];
	assign rdata1 = register_file[raddr1];
	
	//---------------------------------------------------------------
	// Sequential Logic
	//---------------------------------------------------------------
	always @ (posedge clk)
	if (wren) begin
        register_file[waddr]=wdata;
	end
	
	
 endmodule  



